LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY EvenParityChecker IS	
	GENERIC(
	DATAWIDTH: integer:=9
	);
	PORT(
	DATA: IN std_logic_vector(DATAWIDTH-1 DOWNTO 0);
	ENABLE: IN std_logic;
	ERROR: OUT std_logic
	);
END ENTITY EvenParityChecker; 

ARCHITECTURE DataFlow OF EvenParityChecker IS

BEGIN
	
	WITH DATAWIDTH SELECT
	ERROR<=(((((DATA(0) XOR DATA(1)) XOR (DATA(2) XOR DATA(3))) XOR ((DATA(4) XOR DATA(5)) XOR (DATA(6) XOR DATA(7)))) XOR DATA(DATAWIDTH-1))  AND ENABLE)				  
	WHEN 9,(((((DATA(0) XOR DATA(1)) XOR (DATA(2) XOR DATA(3))) XOR ((DATA(4) XOR DATA(5)) XOR (DATA(6) XOR '0'))) XOR DATA(7))  AND ENABLE) WHEN 8,
	'0' WHEN OTHERS;

	
END ARCHITECTURE DataFlow;
